package test_pkg;

    import timer_pkg::*;
    `include "base_test.sv"
    `include "def_val_reg_test.sv"
    `include "R_and_W_value_check.sv"
    `include "reset_on_the_fly_check.sv"
    `include "RW1C_check.sv"
    `include "reserved_register_check.sv"
    `include "count_up_0_nod_interrupt_test.sv"
    `include "count_up_0_d2_interrupt_test.sv"
    `include "count_up_0_d4_interrupt_test.sv"
    `include "count_up_0_d8_interrupt_test.sv"
    `include "count_down_255_nod_interrupt_test.sv"
    `include "count_down_255_d2_interrupt_test.sv"
    `include "count_down_255_d4_interrupt_test.sv"
    `include "count_down_255_d8_interrupt_test.sv"
    `include "count_up_rand_nod_interrupt_test.sv"
    `include "count_up_rand_d2_interrupt_test.sv"        
    `include "count_up_rand_d8_interrupt_test.sv"
    `include "count_up_rand_d4_interrupt_test.sv"
    `include "count_down_rand_nod_interrupt_test.sv"
    `include "count_down_rand_d2_interrupt_test.sv"
    `include "count_down_rand_d4_interrupt_test.sv"
    `include "count_down_rand_d8_interrupt_test.sv"
    `include "count_up_0_then_change_the_counter_at_the_middle_interrupt_test.sv"
    `include "count_up_0_then_change_to_count_down_interrupt_test.sv"
    `include "count_down_255_then_change_the_counter_at_the_middle_interrupt_test.sv"
    `include "count_down_255_then_change_to_count_up_interrupt_test.sv"
    `include "count_up_rand_then_change_to_count_down_interrupt_test.sv"
    `include "count_down_rand_then_change_to_count_up_interrupt_test.sv"
    `include "count_down_with_data_change_divide_at_the_middle_test.sv"
    `include "count_down_with_out_data_change_divide_at_the_middle_test.sv"
    `include "count_up_with_data_change_divide_at_the_middle_test.sv"
    `include "count_up_with_out_data_change_divide_at_the_middle_test.sv"
    `include "count_down_with_data_changes_divide_at_the_middle_then_count_up.sv"
    `include "count_down_with_out_data_changes_divide_at_the_middle_then_count_up.sv"
    `include "count_up_with_data_changes_divide_at_the_middle_then_count_down.sv"
    `include "count_up_with_out_data_changes_divide_at_the_middle_then_count_down.sv"
    `include "count_up_with_rand_divde_then_changes_rand_divide.sv"
    `include "count_up_with_data_rand_divde_then_changes_rand_divide.sv"
    `include "count_down_with_rand_divde_then_changes_rand_divide.sv"
    `include "count_down_with_data_rand_divde_then_changes_rand_divide.sv"
endpackage
